`timescale 1ns / 1ps

module interpolatingFilter_tb;

    // Input signals
    reg clk;
    reg clk_enable;
    reg reset;
    reg signed [15:0] input_data;

    // Output signals
    wire signed [15:0] output_data;
    wire ce_out;
	 integer i;
    // Instantiate the top module
    interpolatingFilter uut (
        .clk(clk),
        .clk_enable(clk_enable),
        .reset(reset),
        .input_data(input_data),
        .output_data(output_data),
        .ce_out(ce_out)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #11350 clk = ~clk;  // Generate a 44.1 kHz clock
    end

    // Test stimuli - chirp signal
    reg signed [16:0] filter_in_data_log_force[0:1035];

    initial begin
        // Initialize inputs
        clk_enable = 1;
        reset = 1;
        input_data = 0;

        // Reset the system
        #100;
        reset = 1;
        #100;
        reset = 0;
        #100;

        // Load test data
		 filter_in_data_log_force[   0] <= 17'h00000;
		 filter_in_data_log_force[   1] <= 17'h08000;
		 filter_in_data_log_force[   2] <= 17'h08000;
		 filter_in_data_log_force[   3] <= 17'h08000;
		 filter_in_data_log_force[   4] <= 17'h00000;
		 filter_in_data_log_force[   5] <= 17'h00000;
		 filter_in_data_log_force[   6] <= 17'h00000;
		 filter_in_data_log_force[   7] <= 17'h00000;				
		 filter_in_data_log_force[   8] <= 17'h08000;
		 filter_in_data_log_force[   9] <= 17'h08000;
		 filter_in_data_log_force[  10] <= 17'h07fff;
		 filter_in_data_log_force[  11] <= 17'h07ffd;
		 filter_in_data_log_force[  12] <= 17'h07ff7;
		 filter_in_data_log_force[  13] <= 17'h07fe9;
		 filter_in_data_log_force[  14] <= 17'h07fd0;
		 filter_in_data_log_force[  15] <= 17'h07fa7;
		 filter_in_data_log_force[  16] <= 17'h07f68;
		 filter_in_data_log_force[  17] <= 17'h07f0d;
		 filter_in_data_log_force[  18] <= 17'h07e8e;
		 filter_in_data_log_force[  19] <= 17'h07de2;
		 filter_in_data_log_force[  20] <= 17'h07d02;
		 filter_in_data_log_force[  21] <= 17'h07be2;
		 filter_in_data_log_force[  22] <= 17'h07a79;
		 filter_in_data_log_force[  23] <= 17'h078bc;
		 filter_in_data_log_force[  24] <= 17'h0769f;
		 filter_in_data_log_force[  25] <= 17'h07416;
		 filter_in_data_log_force[  26] <= 17'h07116;
		 filter_in_data_log_force[  27] <= 17'h06d93;
		 filter_in_data_log_force[  28] <= 17'h06981;
		 filter_in_data_log_force[  29] <= 17'h064d6;
		 filter_in_data_log_force[  30] <= 17'h05f87;
		 filter_in_data_log_force[  31] <= 17'h0598b;
		 filter_in_data_log_force[  32] <= 17'h052db;
		 filter_in_data_log_force[  33] <= 17'h04b71;
		 filter_in_data_log_force[  34] <= 17'h0434b;
		 filter_in_data_log_force[  35] <= 17'h03a68;
		 filter_in_data_log_force[  36] <= 17'h030ca;
		 filter_in_data_log_force[  37] <= 17'h02679;
		 filter_in_data_log_force[  38] <= 17'h01b7f;
		 filter_in_data_log_force[  39] <= 17'h00fec;
		 filter_in_data_log_force[  40] <= 17'h003d4;
		 filter_in_data_log_force[  41] <= 17'h1f751;
		 filter_in_data_log_force[  42] <= 17'h1ea82;
		 filter_in_data_log_force[  43] <= 17'h1dd8b;
		 filter_in_data_log_force[  44] <= 17'h1d098;
		 filter_in_data_log_force[  45] <= 17'h1c3d9;
		 filter_in_data_log_force[  46] <= 17'h1b781;
		 filter_in_data_log_force[  47] <= 17'h1abcc;
		 filter_in_data_log_force[  48] <= 17'h1a0f5;
		 filter_in_data_log_force[  49] <= 17'h1973d;
		 filter_in_data_log_force[  50] <= 17'h18ee4;
		 filter_in_data_log_force[  51] <= 17'h1882c;
		 filter_in_data_log_force[  52] <= 17'h18353;
		 filter_in_data_log_force[  53] <= 17'h18092;
		 filter_in_data_log_force[  54] <= 17'h1801e;
		 filter_in_data_log_force[  55] <= 17'h18220;
		 filter_in_data_log_force[  56] <= 17'h186b8;
		 filter_in_data_log_force[  57] <= 17'h18df5;
		 filter_in_data_log_force[  58] <= 17'h197d9;
		 filter_in_data_log_force[  59] <= 17'h1a450;
		 filter_in_data_log_force[  60] <= 17'h1b334;
		 filter_in_data_log_force[  61] <= 17'h1c445;
		 filter_in_data_log_force[  62] <= 17'h1d731;
		 filter_in_data_log_force[  63] <= 17'h1eb8d;
		 filter_in_data_log_force[  64] <= 17'h000d7;
		 filter_in_data_log_force[  65] <= 17'h0167d;
		 filter_in_data_log_force[  66] <= 17'h02bda;
		 filter_in_data_log_force[  67] <= 17'h0403c;
		 filter_in_data_log_force[  68] <= 17'h052ed;
		 filter_in_data_log_force[  69] <= 17'h06336;
		 filter_in_data_log_force[  70] <= 17'h07067;
		 filter_in_data_log_force[  71] <= 17'h079df;
		 filter_in_data_log_force[  72] <= 17'h07f16;
		 filter_in_data_log_force[  73] <= 17'h07fa5;
		 filter_in_data_log_force[  74] <= 17'h07b4f;
		 filter_in_data_log_force[  75] <= 17'h07205;
		 filter_in_data_log_force[  76] <= 17'h063f1;
		 filter_in_data_log_force[  77] <= 17'h05174;
		 filter_in_data_log_force[  78] <= 17'h03b2d;
		 filter_in_data_log_force[  79] <= 17'h021f3;
		 filter_in_data_log_force[  80] <= 17'h006d0;
		 filter_in_data_log_force[  81] <= 17'h1eafc;
		 filter_in_data_log_force[  82] <= 17'h1cfcb;
		 filter_in_data_log_force[  83] <= 17'h1b6a3;
		 filter_in_data_log_force[  84] <= 17'h1a0e5;
		 filter_in_data_log_force[  85] <= 17'h18fdb;
		 filter_in_data_log_force[  86] <= 17'h184a1;
		 filter_in_data_log_force[  87] <= 17'h18012;
		 filter_in_data_log_force[  88] <= 17'h182b3;
		 filter_in_data_log_force[  89] <= 17'h18ca2;
		 filter_in_data_log_force[  90] <= 17'h19d8d;
		 filter_in_data_log_force[  91] <= 17'h1b4ac;
		 filter_in_data_log_force[  92] <= 17'h1d0c5;
		 filter_in_data_log_force[  93] <= 17'h1f038;
		 filter_in_data_log_force[  94] <= 17'h01110;
		 filter_in_data_log_force[  95] <= 17'h03124;
		 filter_in_data_log_force[  96] <= 17'h04e36;
		 filter_in_data_log_force[  97] <= 17'h06620;
		 filter_in_data_log_force[  98] <= 17'h076fa;
		 filter_in_data_log_force[  99] <= 17'h07f4a;
		 filter_in_data_log_force[ 100] <= 17'h07e28;
		 filter_in_data_log_force[ 101] <= 17'h07359;
		 filter_in_data_log_force[ 102] <= 17'h05f67;
		 filter_in_data_log_force[ 103] <= 17'h043a0;
		 filter_in_data_log_force[ 104] <= 17'h0220b;
		 filter_in_data_log_force[ 105] <= 17'h1fd49;
		 filter_in_data_log_force[ 106] <= 17'h1d863;
		 filter_in_data_log_force[ 107] <= 17'h1b68f;
		 filter_in_data_log_force[ 108] <= 17'h19ae7;
		 filter_in_data_log_force[ 109] <= 17'h1881b;
		 filter_in_data_log_force[ 110] <= 17'h1802d;
		 filter_in_data_log_force[ 111] <= 17'h1842d;
		 filter_in_data_log_force[ 112] <= 17'h19413;
		 filter_in_data_log_force[ 113] <= 17'h1aea8;
		 filter_in_data_log_force[ 114] <= 17'h1d193;
		 filter_in_data_log_force[ 115] <= 17'h1f985;
		 filter_in_data_log_force[ 116] <= 17'h0227f;
		 filter_in_data_log_force[ 117] <= 17'h04837;
		 filter_in_data_log_force[ 118] <= 17'h06687;
		 filter_in_data_log_force[ 119] <= 17'h079ed;
		 filter_in_data_log_force[ 120] <= 17'h07ff5;
		 filter_in_data_log_force[ 121] <= 17'h07793;
		 filter_in_data_log_force[ 122] <= 17'h0615e;
		 filter_in_data_log_force[ 123] <= 17'h03f93;
		 filter_in_data_log_force[ 124] <= 17'h015ed;
		 filter_in_data_log_force[ 125] <= 17'h1e947;
		 filter_in_data_log_force[ 126] <= 17'h1bf10;
		 filter_in_data_log_force[ 127] <= 17'h19ca4;
		 filter_in_data_log_force[ 128] <= 17'h18699;
		 filter_in_data_log_force[ 129] <= 17'h1801a;
		 filter_in_data_log_force[ 130] <= 17'h18a66;
		 filter_in_data_log_force[ 131] <= 17'h1a483;
		 filter_in_data_log_force[ 132] <= 17'h1cb45;
		 filter_in_data_log_force[ 133] <= 17'h1f99d;
		 filter_in_data_log_force[ 134] <= 17'h02936;
		 filter_in_data_log_force[ 135] <= 17'h0534a;
		 filter_in_data_log_force[ 136] <= 17'h0719f;
		 filter_in_data_log_force[ 137] <= 17'h07f76;
		 filter_in_data_log_force[ 138] <= 17'h07a5d;
		 filter_in_data_log_force[ 139] <= 17'h062ab;
		 filter_in_data_log_force[ 140] <= 17'h03b9c;
		 filter_in_data_log_force[ 141] <= 17'h00af3;
		 filter_in_data_log_force[ 142] <= 17'h1d835;
		 filter_in_data_log_force[ 143] <= 17'h1ab83;
		 filter_in_data_log_force[ 144] <= 17'h18c4e;
		 filter_in_data_log_force[ 145] <= 17'h18010;
		 filter_in_data_log_force[ 146] <= 17'h18940;
		 filter_in_data_log_force[ 147] <= 17'h1a6c3;
		 filter_in_data_log_force[ 148] <= 17'h1d3ea;
		 filter_in_data_log_force[ 149] <= 17'h0091c;
		 filter_in_data_log_force[ 150] <= 17'h03d09;
		 filter_in_data_log_force[ 151] <= 17'h0664b;
		 filter_in_data_log_force[ 152] <= 17'h07d1b;
		 filter_in_data_log_force[ 153] <= 17'h07cdd;
		 filter_in_data_log_force[ 154] <= 17'h06523;
		 filter_in_data_log_force[ 155] <= 17'h039fc;
		 filter_in_data_log_force[ 156] <= 17'h0035b;
		 filter_in_data_log_force[ 157] <= 17'h1cbba;
		 filter_in_data_log_force[ 158] <= 17'h19e1d;
		 filter_in_data_log_force[ 159] <= 17'h183e4;
		 filter_in_data_log_force[ 160] <= 17'h182c7;
		 filter_in_data_log_force[ 161] <= 17'h19b7c;
		 filter_in_data_log_force[ 162] <= 17'h1c958;
		 filter_in_data_log_force[ 163] <= 17'h0030c;
		 filter_in_data_log_force[ 164] <= 17'h03c71;
		 filter_in_data_log_force[ 165] <= 17'h0690f;
		 filter_in_data_log_force[ 166] <= 17'h07eda;
		 filter_in_data_log_force[ 167] <= 17'h0788b;
		 filter_in_data_log_force[ 168] <= 17'h0570b;
		 filter_in_data_log_force[ 169] <= 17'h0217e;
		 filter_in_data_log_force[ 170] <= 17'h1e3e8;
		 filter_in_data_log_force[ 171] <= 17'h1ac88;
		 filter_in_data_log_force[ 172] <= 17'h18896;
		 filter_in_data_log_force[ 173] <= 17'h18107;
		 filter_in_data_log_force[ 174] <= 17'h1982e;
		 filter_in_data_log_force[ 175] <= 17'h1c8e8;
		 filter_in_data_log_force[ 176] <= 17'h00791;
		 filter_in_data_log_force[ 177] <= 17'h044ab;
		 filter_in_data_log_force[ 178] <= 17'h070ac;
		 filter_in_data_log_force[ 179] <= 17'h07ffa;
		 filter_in_data_log_force[ 180] <= 17'h06e20;
		 filter_in_data_log_force[ 181] <= 17'h03f3f;
		 filter_in_data_log_force[ 182] <= 17'h1ff51;
		 filter_in_data_log_force[ 183] <= 17'h1bf3c;
		 filter_in_data_log_force[ 184] <= 17'h1906c;
		 filter_in_data_log_force[ 185] <= 17'h18006;
		 filter_in_data_log_force[ 186] <= 17'h19319;
		 filter_in_data_log_force[ 187] <= 17'h1c4db;
		 filter_in_data_log_force[ 188] <= 17'h007a9;
		 filter_in_data_log_force[ 189] <= 17'h0489a;
		 filter_in_data_log_force[ 190] <= 17'h074cd;
		 filter_in_data_log_force[ 191] <= 17'h07ef5;
		 filter_in_data_log_force[ 192] <= 17'h06387;
		 filter_in_data_log_force[ 193] <= 17'h02a25;
		 filter_in_data_log_force[ 194] <= 17'h1e3b9;
		 filter_in_data_log_force[ 195] <= 17'h1a59d;
		 filter_in_data_log_force[ 196] <= 17'h18327;
		 filter_in_data_log_force[ 197] <= 17'h18789;
		 filter_in_data_log_force[ 198] <= 17'h1b1f6;
		 filter_in_data_log_force[ 199] <= 17'h1f579;
		 filter_in_data_log_force[ 200] <= 17'h03cb1;
		 filter_in_data_log_force[ 201] <= 17'h0707c;
		 filter_in_data_log_force[ 202] <= 17'h07f8a;
		 filter_in_data_log_force[ 203] <= 17'h0644f;
		 filter_in_data_log_force[ 204] <= 17'h02751;
		 filter_in_data_log_force[ 205] <= 17'h1dcba;
		 filter_in_data_log_force[ 206] <= 17'h19ddf;
		 filter_in_data_log_force[ 207] <= 17'h180a3;
		 filter_in_data_log_force[ 208] <= 17'h18fb4;
		 filter_in_data_log_force[ 209] <= 17'h1c665;
		 filter_in_data_log_force[ 210] <= 17'h011d0;
		 filter_in_data_log_force[ 211] <= 17'h05729;
		 filter_in_data_log_force[ 212] <= 17'h07d35;
		 filter_in_data_log_force[ 213] <= 17'h07596;
		 filter_in_data_log_force[ 214] <= 17'h0427d;
		 filter_in_data_log_force[ 215] <= 17'h1f660;
		 filter_in_data_log_force[ 216] <= 17'h1ad91;
		 filter_in_data_log_force[ 217] <= 17'h183c7;
		 filter_in_data_log_force[ 218] <= 17'h18977;
		 filter_in_data_log_force[ 219] <= 17'h1bd0f;
		 filter_in_data_log_force[ 220] <= 17'h00b04;
		 filter_in_data_log_force[ 221] <= 17'h054f3;
		 filter_in_data_log_force[ 222] <= 17'h07d62;
		 filter_in_data_log_force[ 223] <= 17'h073a5;
		 filter_in_data_log_force[ 224] <= 17'h03b06;
		 filter_in_data_log_force[ 225] <= 17'h1ea0e;
		 filter_in_data_log_force[ 226] <= 17'h1a1d0;
		 filter_in_data_log_force[ 227] <= 17'h1807a;
		 filter_in_data_log_force[ 228] <= 17'h19488;
		 filter_in_data_log_force[ 229] <= 17'h1d62b;
		 filter_in_data_log_force[ 230] <= 17'h029ed;
		 filter_in_data_log_force[ 231] <= 17'h06bf0;
		 filter_in_data_log_force[ 232] <= 17'h07f4b;
		 filter_in_data_log_force[ 233] <= 17'h05aed;
		 filter_in_data_log_force[ 234] <= 17'h00e39;
		 filter_in_data_log_force[ 235] <= 17'h1bae5;
		 filter_in_data_log_force[ 236] <= 17'h18655;
		 filter_in_data_log_force[ 237] <= 17'h188c0;
		 filter_in_data_log_force[ 238] <= 17'h1c1b6;
		 filter_in_data_log_force[ 239] <= 17'h0179a;
		 filter_in_data_log_force[ 240] <= 17'h062d5;
		 filter_in_data_log_force[ 241] <= 17'h07ffe;
		 filter_in_data_log_force[ 242] <= 17'h060c0;
		 filter_in_data_log_force[ 243] <= 17'h01349;
		 filter_in_data_log_force[ 244] <= 17'h1bc47;
		 filter_in_data_log_force[ 245] <= 17'h185c6;
		 filter_in_data_log_force[ 246] <= 17'h18ac6;
		 filter_in_data_log_force[ 247] <= 17'h1c981;
		 filter_in_data_log_force[ 248] <= 17'h0237f;
		 filter_in_data_log_force[ 249] <= 17'h06c0a;
		 filter_in_data_log_force[ 250] <= 17'h07e59;
		 filter_in_data_log_force[ 251] <= 17'h05081;
		 filter_in_data_log_force[ 252] <= 17'h1f944;
		 filter_in_data_log_force[ 253] <= 17'h1a536;
		 filter_in_data_log_force[ 254] <= 17'h1801f;
		 filter_in_data_log_force[ 255] <= 17'h19df7;
		 filter_in_data_log_force[ 256] <= 17'h1efb7;
		 filter_in_data_log_force[ 257] <= 17'h04a67;
		 filter_in_data_log_force[ 258] <= 17'h07d75;
		 filter_in_data_log_force[ 259] <= 17'h06cd6;
		 filter_in_data_log_force[ 260] <= 17'h020dc;
		 filter_in_data_log_force[ 261] <= 17'h1c29a;
		 filter_in_data_log_force[ 262] <= 17'h18602;
		 filter_in_data_log_force[ 263] <= 17'h18d36;
		 filter_in_data_log_force[ 264] <= 17'h1d4e4;
		 filter_in_data_log_force[ 265] <= 17'h0352d;
		 filter_in_data_log_force[ 266] <= 17'h07775;
		 filter_in_data_log_force[ 267] <= 17'h0755d;
		 filter_in_data_log_force[ 268] <= 17'h02f64;
		 filter_in_data_log_force[ 269] <= 17'h1cd99;
		 filter_in_data_log_force[ 270] <= 17'h18916;
		 filter_in_data_log_force[ 271] <= 17'h18aa8;
		 filter_in_data_log_force[ 272] <= 17'h1d217;
		 filter_in_data_log_force[ 273] <= 17'h03543;
		 filter_in_data_log_force[ 274] <= 17'h07890;
		 filter_in_data_log_force[ 275] <= 17'h072ba;
		 filter_in_data_log_force[ 276] <= 17'h02699;
		 filter_in_data_log_force[ 277] <= 17'h1c26f;
		 filter_in_data_log_force[ 278] <= 17'h1843c;
		 filter_in_data_log_force[ 279] <= 17'h1934a;
		 filter_in_data_log_force[ 280] <= 17'h1e6e0;
		 filter_in_data_log_force[ 281] <= 17'h04aa2;
		 filter_in_data_log_force[ 282] <= 17'h07f00;
		 filter_in_data_log_force[ 283] <= 17'h061d2;
		 filter_in_data_log_force[ 284] <= 17'h00536;
		 filter_in_data_log_force[ 285] <= 17'h1a4f2;
		 filter_in_data_log_force[ 286] <= 17'h18033;
		 filter_in_data_log_force[ 287] <= 17'h1afd4;
		 filter_in_data_log_force[ 288] <= 17'h014ef;
		 filter_in_data_log_force[ 289] <= 17'h06c4a;
		 filter_in_data_log_force[ 290] <= 17'h07ad7;
		 filter_in_data_log_force[ 291] <= 17'h03607;
		 filter_in_data_log_force[ 292] <= 17'h1cc1a;
		 filter_in_data_log_force[ 293] <= 17'h1859c;
		 filter_in_data_log_force[ 294] <= 17'h193b2;
		 filter_in_data_log_force[ 295] <= 17'h1ed52;
		 filter_in_data_log_force[ 296] <= 17'h05449;
		 filter_in_data_log_force[ 297] <= 17'h07ffc;
		 filter_in_data_log_force[ 298] <= 17'h050d0;
		 filter_in_data_log_force[ 299] <= 17'h1e7b4;
		 filter_in_data_log_force[ 300] <= 17'h18fd3;
		 filter_in_data_log_force[ 301] <= 17'h18906;
		 filter_in_data_log_force[ 302] <= 17'h1d8fc;
		 filter_in_data_log_force[ 303] <= 17'h045c8;
		 filter_in_data_log_force[ 304] <= 17'h07f4c;
		 filter_in_data_log_force[ 305] <= 17'h05a53;
		 filter_in_data_log_force[ 306] <= 17'h1f1b3;
		 filter_in_data_log_force[ 307] <= 17'h19396;
		 filter_in_data_log_force[ 308] <= 17'h1875d;
		 filter_in_data_log_force[ 309] <= 17'h1d710;
		 filter_in_data_log_force[ 310] <= 17'h04658;
		 filter_in_data_log_force[ 311] <= 17'h07f9b;
		 filter_in_data_log_force[ 312] <= 17'h055ee;
		 filter_in_data_log_force[ 313] <= 17'h1e908;
		 filter_in_data_log_force[ 314] <= 17'h18def;
		 filter_in_data_log_force[ 315] <= 17'h18cd3;
		 filter_in_data_log_force[ 316] <= 17'h1e756;
		 filter_in_data_log_force[ 317] <= 17'h055cb;
		 filter_in_data_log_force[ 318] <= 17'h07f6c;
		 filter_in_data_log_force[ 319] <= 17'h041ef;
		 filter_in_data_log_force[ 320] <= 17'h1ce96;
		 filter_in_data_log_force[ 321] <= 17'h1837d;
		 filter_in_data_log_force[ 322] <= 17'h19ee4;
		 filter_in_data_log_force[ 323] <= 17'h00ae5;
		 filter_in_data_log_force[ 324] <= 17'h06e0b;
		 filter_in_data_log_force[ 325] <= 17'h0750f;
		 filter_in_data_log_force[ 326] <= 17'h01948;
		 filter_in_data_log_force[ 327] <= 17'h1a7d8;
		 filter_in_data_log_force[ 328] <= 17'h18172;
		 filter_in_data_log_force[ 329] <= 17'h1c7a9;
		 filter_in_data_log_force[ 330] <= 17'h03eb0;
		 filter_in_data_log_force[ 331] <= 17'h07f80;
		 filter_in_data_log_force[ 332] <= 17'h0510b;
		 filter_in_data_log_force[ 333] <= 17'h1db47;
		 filter_in_data_log_force[ 334] <= 17'h185ba;
		 filter_in_data_log_force[ 335] <= 17'h19caa;
		 filter_in_data_log_force[ 336] <= 17'h00c6d;
		 filter_in_data_log_force[ 337] <= 17'h0713e;
		 filter_in_data_log_force[ 338] <= 17'h06feb;
		 filter_in_data_log_force[ 339] <= 17'h008e1;
		 filter_in_data_log_force[ 340] <= 17'h19987;
		 filter_in_data_log_force[ 341] <= 17'h1881f;
		 filter_in_data_log_force[ 342] <= 17'h1e571;
		 filter_in_data_log_force[ 343] <= 17'h05b9d;
		 filter_in_data_log_force[ 344] <= 17'h07c6f;
		 filter_in_data_log_force[ 345] <= 17'h02872;
		 filter_in_data_log_force[ 346] <= 17'h1ae1b;
		 filter_in_data_log_force[ 347] <= 17'h1814b;
		 filter_in_data_log_force[ 348] <= 17'h1cd58;
		 filter_in_data_log_force[ 349] <= 17'h04a26;
		 filter_in_data_log_force[ 350] <= 17'h07fa4;
		 filter_in_data_log_force[ 351] <= 17'h0396c;
		 filter_in_data_log_force[ 352] <= 17'h1bb15;
		 filter_in_data_log_force[ 353] <= 17'h18014;
		 filter_in_data_log_force[ 354] <= 17'h1c308;
		 filter_in_data_log_force[ 355] <= 17'h04281;
		 filter_in_data_log_force[ 356] <= 17'h07ff9;
		 filter_in_data_log_force[ 357] <= 17'h03d6f;
		 filter_in_data_log_force[ 358] <= 17'h1bcf6;
		 filter_in_data_log_force[ 359] <= 17'h18014;
		 filter_in_data_log_force[ 360] <= 17'h1c529;
		 filter_in_data_log_force[ 361] <= 17'h0467d;
		 filter_in_data_log_force[ 362] <= 17'h07fa1;
		 filter_in_data_log_force[ 363] <= 17'h03515;
		 filter_in_data_log_force[ 364] <= 17'h1b354;
		 filter_in_data_log_force[ 365] <= 17'h18155;
		 filter_in_data_log_force[ 366] <= 17'h1d40c;
		 filter_in_data_log_force[ 367] <= 17'h05535;
		 filter_in_data_log_force[ 368] <= 17'h07c58;
		 filter_in_data_log_force[ 369] <= 17'h01f36;
		 filter_in_data_log_force[ 370] <= 17'h1a08c;
		 filter_in_data_log_force[ 371] <= 17'h18849;
		 filter_in_data_log_force[ 372] <= 17'h1f14f;
		 filter_in_data_log_force[ 373] <= 17'h06a71;
		 filter_in_data_log_force[ 374] <= 17'h06fa4;
		 filter_in_data_log_force[ 375] <= 17'h1fa75;
		 filter_in_data_log_force[ 376] <= 17'h18b33;
		 filter_in_data_log_force[ 377] <= 17'h19d15;
		 filter_in_data_log_force[ 378] <= 17'h01d08;
		 filter_in_data_log_force[ 379] <= 17'h07cb8;
		 filter_in_data_log_force[ 380] <= 17'h05075;
		 filter_in_data_log_force[ 381] <= 17'h1c953;
		 filter_in_data_log_force[ 382] <= 17'h18000;
		 filter_in_data_log_force[ 383] <= 17'h1c86d;
		 filter_in_data_log_force[ 384] <= 17'h05095;
		 filter_in_data_log_force[ 385] <= 17'h07c3b;
		 filter_in_data_log_force[ 386] <= 17'h0185b;
		 filter_in_data_log_force[ 387] <= 17'h1980f;
		 filter_in_data_log_force[ 388] <= 17'h190db;
		 filter_in_data_log_force[ 389] <= 17'h00bee;
		 filter_in_data_log_force[ 390] <= 17'h0791f;
		 filter_in_data_log_force[ 391] <= 17'h05727;
		 filter_in_data_log_force[ 392] <= 17'h1cd8b;
		 filter_in_data_log_force[ 393] <= 17'h18001;
		 filter_in_data_log_force[ 394] <= 17'h1cbeb;
		 filter_in_data_log_force[ 395] <= 17'h056b3;
		 filter_in_data_log_force[ 396] <= 17'h078b1;
		 filter_in_data_log_force[ 397] <= 17'h007f0;
		 filter_in_data_log_force[ 398] <= 17'h18d58;
		 filter_in_data_log_force[ 399] <= 17'h19f50;
		 filter_in_data_log_force[ 400] <= 17'h02883;
		 filter_in_data_log_force[ 401] <= 17'h07fb5;
		 filter_in_data_log_force[ 402] <= 17'h03825;
		 filter_in_data_log_force[ 403] <= 17'h1aa56;
		 filter_in_data_log_force[ 404] <= 17'h187e1;
		 filter_in_data_log_force[ 405] <= 17'h1fcd2;
		 filter_in_data_log_force[ 406] <= 17'h075ee;
		 filter_in_data_log_force[ 407] <= 17'h0592f;
		 filter_in_data_log_force[ 408] <= 17'h1ca78;
		 filter_in_data_log_force[ 409] <= 17'h18047;
		 filter_in_data_log_force[ 410] <= 17'h1da9b;
		 filter_in_data_log_force[ 411] <= 17'h06570;
		 filter_in_data_log_force[ 412] <= 17'h06c8e;
		 filter_in_data_log_force[ 413] <= 17'h1e5f2;
		 filter_in_data_log_force[ 414] <= 17'h1815a;
		 filter_in_data_log_force[ 415] <= 17'h1c370;
		 filter_in_data_log_force[ 416] <= 17'h055b2;
		 filter_in_data_log_force[ 417] <= 17'h07649;
		 filter_in_data_log_force[ 418] <= 17'h1f920;
		 filter_in_data_log_force[ 419] <= 17'h1850b;
		 filter_in_data_log_force[ 420] <= 17'h1b641;
		 filter_in_data_log_force[ 421] <= 17'h04b25;
		 filter_in_data_log_force[ 422] <= 17'h07a3e;
		 filter_in_data_log_force[ 423] <= 17'h002da;
		 filter_in_data_log_force[ 424] <= 17'h18770;
		 filter_in_data_log_force[ 425] <= 17'h1b187;
		 filter_in_data_log_force[ 426] <= 17'h047e9;
		 filter_in_data_log_force[ 427] <= 17'h07ad4;
		 filter_in_data_log_force[ 428] <= 17'h002f3;
		 filter_in_data_log_force[ 429] <= 17'h186d6;
		 filter_in_data_log_force[ 430] <= 17'h1b487;
		 filter_in_data_log_force[ 431] <= 17'h04c8a;
		 filter_in_data_log_force[ 432] <= 17'h07879;
		 filter_in_data_log_force[ 433] <= 17'h1f96b;
		 filter_in_data_log_force[ 434] <= 17'h183a2;
		 filter_in_data_log_force[ 435] <= 17'h1bfbb;
		 filter_in_data_log_force[ 436] <= 17'h0583c;
		 filter_in_data_log_force[ 437] <= 17'h07193;
		 filter_in_data_log_force[ 438] <= 17'h1e66d;
		 filter_in_data_log_force[ 439] <= 17'h1805a;
		 filter_in_data_log_force[ 440] <= 17'h1d490;
		 filter_in_data_log_force[ 441] <= 17'h06885;
		 filter_in_data_log_force[ 442] <= 17'h062c8;
		 filter_in_data_log_force[ 443] <= 17'h1cb18;
		 filter_in_data_log_force[ 444] <= 17'h181c2;
		 filter_in_data_log_force[ 445] <= 17'h1f458;
		 filter_in_data_log_force[ 446] <= 17'h07872;
		 filter_in_data_log_force[ 447] <= 17'h047e5;
		 filter_in_data_log_force[ 448] <= 17'h1aaff;
		 filter_in_data_log_force[ 449] <= 17'h18e89;
		 filter_in_data_log_force[ 450] <= 17'h01e51;
		 filter_in_data_log_force[ 451] <= 17'h08000;
		 filter_in_data_log_force[ 452] <= 17'h01def;
		 filter_in_data_log_force[ 453] <= 17'h18dd4;
		 filter_in_data_log_force[ 454] <= 17'h1ada0;
		 filter_in_data_log_force[ 455] <= 17'h04cea;
		 filter_in_data_log_force[ 456] <= 17'h074d8;
		 filter_in_data_log_force[ 457] <= 17'h1e69f;
		 filter_in_data_log_force[ 458] <= 17'h18006;
		 filter_in_data_log_force[ 459] <= 17'h1e264;
		 filter_in_data_log_force[ 460] <= 17'h07383;
		 filter_in_data_log_force[ 461] <= 17'h04de9;
		 filter_in_data_log_force[ 462] <= 17'h1ac86;
		 filter_in_data_log_force[ 463] <= 17'h19022;
		 filter_in_data_log_force[ 464] <= 17'h026bf;
		 filter_in_data_log_force[ 465] <= 17'h07f38;
		 filter_in_data_log_force[ 466] <= 17'h00aa8;
		 filter_in_data_log_force[ 467] <= 17'h184c9;
		 filter_in_data_log_force[ 468] <= 17'h1c6ed;
		 filter_in_data_log_force[ 469] <= 17'h06620;
		 filter_in_data_log_force[ 470] <= 17'h05e5e;
		 filter_in_data_log_force[ 471] <= 17'h1bbb1;
		 filter_in_data_log_force[ 472] <= 17'h18978;
		 filter_in_data_log_force[ 473] <= 17'h01b35;
		 filter_in_data_log_force[ 474] <= 17'h07fe0;
		 filter_in_data_log_force[ 475] <= 17'h00fa4;
		 filter_in_data_log_force[ 476] <= 17'h18536;
		 filter_in_data_log_force[ 477] <= 17'h1c8a7;
		 filter_in_data_log_force[ 478] <= 17'h06948;
		 filter_in_data_log_force[ 479] <= 17'h0582a;
		 filter_in_data_log_force[ 480] <= 17'h1b19a;
		 filter_in_data_log_force[ 481] <= 17'h19051;
		 filter_in_data_log_force[ 482] <= 17'h02da6;
		 filter_in_data_log_force[ 483] <= 17'h07cdd;
		 filter_in_data_log_force[ 484] <= 17'h1f580;
		 filter_in_data_log_force[ 485] <= 17'h18031;
		 filter_in_data_log_force[ 486] <= 17'h1e808;
		 filter_in_data_log_force[ 487] <= 17'h0798a;
		 filter_in_data_log_force[ 488] <= 17'h0374f;
		 filter_in_data_log_force[ 489] <= 17'h19458;
		 filter_in_data_log_force[ 490] <= 17'h1ae34;
		 filter_in_data_log_force[ 491] <= 17'h05814;
		 filter_in_data_log_force[ 492] <= 17'h0666d;
		 filter_in_data_log_force[ 493] <= 17'h1bf3c;
		 filter_in_data_log_force[ 494] <= 17'h18b2b;
		 filter_in_data_log_force[ 495] <= 17'h0278f;
		 filter_in_data_log_force[ 496] <= 17'h07d2c;
		 filter_in_data_log_force[ 497] <= 17'h1f1f6;
		 filter_in_data_log_force[ 498] <= 17'h18002;
		 filter_in_data_log_force[ 499] <= 17'h1f579;
		 filter_in_data_log_force[ 500] <= 17'h07e12;
		 filter_in_data_log_force[ 501] <= 17'h02138;
		 filter_in_data_log_force[ 502] <= 17'h187ae;
		 filter_in_data_log_force[ 503] <= 17'h1ca8f;
		 filter_in_data_log_force[ 504] <= 17'h06fb2;
		 filter_in_data_log_force[ 505] <= 17'h046e0;
		 filter_in_data_log_force[ 506] <= 17'h19ae9;
		 filter_in_data_log_force[ 507] <= 17'h1aa8e;
		 filter_in_data_log_force[ 508] <= 17'h05952;
		 filter_in_data_log_force[ 509] <= 17'h06140;
		 filter_in_data_log_force[ 510] <= 17'h1b2ea;
		 filter_in_data_log_force[ 511] <= 17'h1957c;
		 filter_in_data_log_force[ 512] <= 17'h040f7;
		 filter_in_data_log_force[ 513] <= 17'h0718c;
		 filter_in_data_log_force[ 514] <= 17'h1ca99;
		 filter_in_data_log_force[ 515] <= 17'h18951;
		 filter_in_data_log_force[ 516] <= 17'h02abe;
		 filter_in_data_log_force[ 517] <= 17'h07a48;
		 filter_in_data_log_force[ 518] <= 17'h1dec7;
		 filter_in_data_log_force[ 519] <= 17'h18351;
		 filter_in_data_log_force[ 520] <= 17'h01905;
		 filter_in_data_log_force[ 521] <= 17'h07e31;
		 filter_in_data_log_force[ 522] <= 17'h1edc5;
		 filter_in_data_log_force[ 523] <= 17'h180ee;
		 filter_in_data_log_force[ 524] <= 17'h00ced;
		 filter_in_data_log_force[ 525] <= 17'h07f8a;
		 filter_in_data_log_force[ 526] <= 17'h1f6dd;
		 filter_in_data_log_force[ 527] <= 17'h1803d;
		 filter_in_data_log_force[ 528] <= 17'h006e0;
		 filter_in_data_log_force[ 529] <= 17'h07fd8;
		 filter_in_data_log_force[ 530] <= 17'h1f9d9;
		 filter_in_data_log_force[ 531] <= 17'h18029;
		 filter_in_data_log_force[ 532] <= 17'h006f8;
		 filter_in_data_log_force[ 533] <= 17'h07fc1;
		 filter_in_data_log_force[ 534] <= 17'h1f6ad;
		 filter_in_data_log_force[ 535] <= 17'h1807b;
		 filter_in_data_log_force[ 536] <= 17'h00d35;
		 filter_in_data_log_force[ 537] <= 17'h07f08;
		 filter_in_data_log_force[ 538] <= 17'h1ed65;
		 filter_in_data_log_force[ 539] <= 17'h181e1;
		 filter_in_data_log_force[ 540] <= 17'h0197b;
		 filter_in_data_log_force[ 541] <= 17'h07c91;
		 filter_in_data_log_force[ 542] <= 17'h1de3b;
		 filter_in_data_log_force[ 543] <= 17'h185e6;
		 filter_in_data_log_force[ 544] <= 17'h02b5d;
		 filter_in_data_log_force[ 545] <= 17'h0766b;
		 filter_in_data_log_force[ 546] <= 17'h1c9ea;
		 filter_in_data_log_force[ 547] <= 17'h18ed4;
		 filter_in_data_log_force[ 548] <= 17'h041b2;
		 filter_in_data_log_force[ 549] <= 17'h06a04;
		 filter_in_data_log_force[ 550] <= 17'h1b229;
		 filter_in_data_log_force[ 551] <= 17'h19f65;
		 filter_in_data_log_force[ 552] <= 17'h05a10;
		 filter_in_data_log_force[ 553] <= 17'h054a3;
		 filter_in_data_log_force[ 554] <= 17'h19a38;
		 filter_in_data_log_force[ 555] <= 17'h1ba1c;
		 filter_in_data_log_force[ 556] <= 17'h0704a;
		 filter_in_data_log_force[ 557] <= 17'h03448;
		 filter_in_data_log_force[ 558] <= 17'h1873c;
		 filter_in_data_log_force[ 559] <= 17'h1e01a;
		 filter_in_data_log_force[ 560] <= 17'h07e4e;
		 filter_in_data_log_force[ 561] <= 17'h00912;
		 filter_in_data_log_force[ 562] <= 17'h18009;
		 filter_in_data_log_force[ 563] <= 17'h00f96;
		 filter_in_data_log_force[ 564] <= 17'h07cd4;
		 filter_in_data_log_force[ 565] <= 17'h1d6e0;
		 filter_in_data_log_force[ 566] <= 17'h18bdf;
		 filter_in_data_log_force[ 567] <= 17'h04244;
		 filter_in_data_log_force[ 568] <= 17'h06557;
		 filter_in_data_log_force[ 569] <= 17'h1a699;
		 filter_in_data_log_force[ 570] <= 17'h1afaa;
		 filter_in_data_log_force[ 571] <= 17'h06cb1;
		 filter_in_data_log_force[ 572] <= 17'h03584;
		 filter_in_data_log_force[ 573] <= 17'h185d7;
		 filter_in_data_log_force[ 574] <= 17'h1ea13;
		 filter_in_data_log_force[ 575] <= 17'h07fe8;
		 filter_in_data_log_force[ 576] <= 17'h1f357;
		 filter_in_data_log_force[ 577] <= 17'h183a5;
		 filter_in_data_log_force[ 578] <= 17'h02fc1;
		 filter_in_data_log_force[ 579] <= 17'h06e8a;
		 filter_in_data_log_force[ 580] <= 17'h1afc0;
		 filter_in_data_log_force[ 581] <= 17'h1a999;
		 filter_in_data_log_force[ 582] <= 17'h06aa8;
		 filter_in_data_log_force[ 583] <= 17'h03515;
		 filter_in_data_log_force[ 584] <= 17'h18484;
		 filter_in_data_log_force[ 585] <= 17'h1f2f0;
		 filter_in_data_log_force[ 586] <= 17'h07fbb;
		 filter_in_data_log_force[ 587] <= 17'h1e22c;
		 filter_in_data_log_force[ 588] <= 17'h18a87;
		 filter_in_data_log_force[ 589] <= 17'h046a6;
		 filter_in_data_log_force[ 590] <= 17'h05c6e;
		 filter_in_data_log_force[ 591] <= 17'h1982b;
		 filter_in_data_log_force[ 592] <= 17'h1c98f;
		 filter_in_data_log_force[ 593] <= 17'h07bfd;
		 filter_in_data_log_force[ 594] <= 17'h007a5;
		 filter_in_data_log_force[ 595] <= 17'h18128;
		 filter_in_data_log_force[ 596] <= 17'h029b4;
		 filter_in_data_log_force[ 597] <= 17'h06e4d;
		 filter_in_data_log_force[ 598] <= 17'h1aa1e;
		 filter_in_data_log_force[ 599] <= 17'h1b4b2;
		 filter_in_data_log_force[ 600] <= 17'h074e5;
		 filter_in_data_log_force[ 601] <= 17'h01a57;
		 filter_in_data_log_force[ 602] <= 17'h18001;
		 filter_in_data_log_force[ 603] <= 17'h01cbe;
		 filter_in_data_log_force[ 604] <= 17'h07360;
		 filter_in_data_log_force[ 605] <= 17'h1b049;
		 filter_in_data_log_force[ 606] <= 17'h1b067;
		 filter_in_data_log_force[ 607] <= 17'h073c5;
		 filter_in_data_log_force[ 608] <= 17'h01a58;
		 filter_in_data_log_force[ 609] <= 17'h1800e;
		 filter_in_data_log_force[ 610] <= 17'h021f8;
		 filter_in_data_log_force[ 611] <= 17'h06fa5;
		 filter_in_data_log_force[ 612] <= 17'h1a825;
		 filter_in_data_log_force[ 613] <= 17'h1bb61;
		 filter_in_data_log_force[ 614] <= 17'h079ba;
		 filter_in_data_log_force[ 615] <= 17'h007a8;
		 filter_in_data_log_force[ 616] <= 17'h1827e;
		 filter_in_data_log_force[ 617] <= 17'h0389d;
		 filter_in_data_log_force[ 618] <= 17'h06017;
		 filter_in_data_log_force[ 619] <= 17'h1951d;
		 filter_in_data_log_force[ 620] <= 17'h1d895;
		 filter_in_data_log_force[ 621] <= 17'h07fe5;
		 filter_in_data_log_force[ 622] <= 17'h1e231;
		 filter_in_data_log_force[ 623] <= 17'h19084;
		 filter_in_data_log_force[ 624] <= 17'h05b64;
		 filter_in_data_log_force[ 625] <= 17'h03c5b;
		 filter_in_data_log_force[ 626] <= 17'h182a4;
		 filter_in_data_log_force[ 627] <= 17'h00b25;
		 filter_in_data_log_force[ 628] <= 17'h076d5;
		 filter_in_data_log_force[ 629] <= 17'h1afc5;
		 filter_in_data_log_force[ 630] <= 17'h1b863;
		 filter_in_data_log_force[ 631] <= 17'h07a9d;
		 filter_in_data_log_force[ 632] <= 17'h1fe23;
		 filter_in_data_log_force[ 633] <= 17'h186a1;
		 filter_in_data_log_force[ 634] <= 17'h04bea;
		 filter_in_data_log_force[ 635] <= 17'h04a80;
		 filter_in_data_log_force[ 636] <= 17'h185da;
		 filter_in_data_log_force[ 637] <= 17'h00232;
		 filter_in_data_log_force[ 638] <= 17'h078a3;
		 filter_in_data_log_force[ 639] <= 17'h1b0c1;
		 filter_in_data_log_force[ 640] <= 17'h1ba8e;
		 filter_in_data_log_force[ 641] <= 17'h07c4f;
		 filter_in_data_log_force[ 642] <= 17'h1f3db;
		 filter_in_data_log_force[ 643] <= 17'h18bdb;
		 filter_in_data_log_force[ 644] <= 17'h0599d;
		 filter_in_data_log_force[ 645] <= 17'h037bb;
		 filter_in_data_log_force[ 646] <= 17'h180ad;
		 filter_in_data_log_force[ 647] <= 17'h01f6f;
		 filter_in_data_log_force[ 648] <= 17'h06981;
		 filter_in_data_log_force[ 649] <= 17'h1973d;
		 filter_in_data_log_force[ 650] <= 17'h1e00e;
		 filter_in_data_log_force[ 651] <= 17'h07f38;
		 filter_in_data_log_force[ 652] <= 17'h1c54c;
		 filter_in_data_log_force[ 653] <= 17'h1ab12;
		 filter_in_data_log_force[ 654] <= 17'h07814;
		 filter_in_data_log_force[ 655] <= 17'h1fd49;
		 filter_in_data_log_force[ 656] <= 17'h18a0f;
		 filter_in_data_log_force[ 657] <= 17'h05a05;
		 filter_in_data_log_force[ 658] <= 17'h032a8;
		 filter_in_data_log_force[ 659] <= 17'h18007;
		 filter_in_data_log_force[ 660] <= 17'h02e47;
		 filter_in_data_log_force[ 661] <= 17'h05c87;
		 filter_in_data_log_force[ 662] <= 17'h18ab6;
		 filter_in_data_log_force[ 663] <= 17'h1fe54;
		 filter_in_data_log_force[ 664] <= 17'h07671;
		 filter_in_data_log_force[ 665] <= 17'h1a4ba;
		 filter_in_data_log_force[ 666] <= 17'h1d1d7;
		 filter_in_data_log_force[ 667] <= 17'h07fe3;
		 filter_in_data_log_force[ 668] <= 17'h1c7a1;
		 filter_in_data_log_force[ 669] <= 17'h1adc3;
		 filter_in_data_log_force[ 670] <= 17'h07b18;
		 filter_in_data_log_force[ 671] <= 17'h1ed78;
		 filter_in_data_log_force[ 672] <= 17'h19454;
		 filter_in_data_log_force[ 673] <= 17'h06bbc;
		 filter_in_data_log_force[ 674] <= 17'h011a8;
		 filter_in_data_log_force[ 675] <= 17'h18598;
		 filter_in_data_log_force[ 676] <= 17'h055d0;
		 filter_in_data_log_force[ 677] <= 17'h03140;
		 filter_in_data_log_force[ 678] <= 17'h18028;
		 filter_in_data_log_force[ 679] <= 17'h03cf1;
		 filter_in_data_log_force[ 680] <= 17'h04ad6;
		 filter_in_data_log_force[ 681] <= 17'h181e0;
		 filter_in_data_log_force[ 682] <= 17'h023f7;
		 filter_in_data_log_force[ 683] <= 17'h05e2f;
		 filter_in_data_log_force[ 684] <= 17'h1886b;
		 filter_in_data_log_force[ 685] <= 17'h00cd6;
		 filter_in_data_log_force[ 686] <= 17'h06bdc;
		 filter_in_data_log_force[ 687] <= 17'h191a0;
		 filter_in_data_log_force[ 688] <= 17'h1f8bb;
		 filter_in_data_log_force[ 689] <= 17'h074db;
		 filter_in_data_log_force[ 690] <= 17'h19bb0;
		 filter_in_data_log_force[ 691] <= 17'h1e834;
		 filter_in_data_log_force[ 692] <= 17'h07a50;
		 filter_in_data_log_force[ 693] <= 17'h1a536;
		 filter_in_data_log_force[ 694] <= 17'h1db63;
		 filter_in_data_log_force[ 695] <= 17'h07d51;
		 filter_in_data_log_force[ 696] <= 17'h1ad34;
		 filter_in_data_log_force[ 697] <= 17'h1d22e;
		 filter_in_data_log_force[ 698] <= 17'h07ec8;
		 filter_in_data_log_force[ 699] <= 17'h1b2ff;
		 filter_in_data_log_force[ 700] <= 17'h1cc64;
		 filter_in_data_log_force[ 701] <= 17'h07f62;
		 filter_in_data_log_force[ 702] <= 17'h1b630;
		 filter_in_data_log_force[ 703] <= 17'h1c9d8;
		 filter_in_data_log_force[ 704] <= 17'h07f88;
		 filter_in_data_log_force[ 705] <= 17'h1b696;
		 filter_in_data_log_force[ 706] <= 17'h1ca75;
		 filter_in_data_log_force[ 707] <= 17'h07f5d;
		 filter_in_data_log_force[ 708] <= 17'h1b429;
		 filter_in_data_log_force[ 709] <= 17'h1ce3e;
		 filter_in_data_log_force[ 710] <= 17'h07eba;
		 filter_in_data_log_force[ 711] <= 17'h1af10;
		 filter_in_data_log_force[ 712] <= 17'h1d555;
		 filter_in_data_log_force[ 713] <= 17'h07d33;
		 filter_in_data_log_force[ 714] <= 17'h1a7a1;
		 filter_in_data_log_force[ 715] <= 17'h1dfec;
		 filter_in_data_log_force[ 716] <= 17'h07a16;
		 filter_in_data_log_force[ 717] <= 17'h19e73;
		 filter_in_data_log_force[ 718] <= 17'h1ee2c;
		 filter_in_data_log_force[ 719] <= 17'h07478;
		 filter_in_data_log_force[ 720] <= 17'h1946a;
		 filter_in_data_log_force[ 721] <= 17'h0001f;
		 filter_in_data_log_force[ 722] <= 17'h06b3f;
		 filter_in_data_log_force[ 723] <= 17'h18ace;
		 filter_in_data_log_force[ 724] <= 17'h0157e;
		 filter_in_data_log_force[ 725] <= 17'h05d49;
		 filter_in_data_log_force[ 726] <= 17'h18350;
		 filter_in_data_log_force[ 727] <= 17'h02d85;
		 filter_in_data_log_force[ 728] <= 17'h0499b;
		 filter_in_data_log_force[ 729] <= 17'h18004;
		 filter_in_data_log_force[ 730] <= 17'h046bc;
		 filter_in_data_log_force[ 731] <= 17'h02fae;
		 filter_in_data_log_force[ 732] <= 17'h18339;
		 filter_in_data_log_force[ 733] <= 17'h05ed9;
		 filter_in_data_log_force[ 734] <= 17'h00fc9;
		 filter_in_data_log_force[ 735] <= 17'h18f2f;
		 filter_in_data_log_force[ 736] <= 17'h072b0;
		 filter_in_data_log_force[ 737] <= 17'h1eb6b;
		 filter_in_data_log_force[ 738] <= 17'h1a58f;
		 filter_in_data_log_force[ 739] <= 17'h07e6d;
		 filter_in_data_log_force[ 740] <= 17'h1c59b;
		 filter_in_data_log_force[ 741] <= 17'h1c6ca;
		 filter_in_data_log_force[ 742] <= 17'h07e15;
		 filter_in_data_log_force[ 743] <= 17'h1a306;
		 filter_in_data_log_force[ 744] <= 17'h1f14f;
		 filter_in_data_log_force[ 745] <= 17'h06e65;
		 filter_in_data_log_force[ 746] <= 17'h189ae;
		 filter_in_data_log_force[ 747] <= 17'h020f4;
		 filter_in_data_log_force[ 748] <= 17'h04e0a;
		 filter_in_data_log_force[ 749] <= 17'h18000;
		 filter_in_data_log_force[ 750] <= 17'h04ec6;
		 filter_in_data_log_force[ 751] <= 17'h01ef0;
		 filter_in_data_log_force[ 752] <= 17'h18b44;
		 filter_in_data_log_force[ 753] <= 17'h071a3;
		 filter_in_data_log_force[ 754] <= 17'h1e742;
		 filter_in_data_log_force[ 755] <= 17'h1ad7f;
		 filter_in_data_log_force[ 756] <= 17'h07ff8;
		 filter_in_data_log_force[ 757] <= 17'h1b180;
		 filter_in_data_log_force[ 758] <= 17'h1e35a;
		 filter_in_data_log_force[ 759] <= 17'h07293;
		 filter_in_data_log_force[ 760] <= 17'h18b02;
		 filter_in_data_log_force[ 761] <= 17'h022e5;
		 filter_in_data_log_force[ 762] <= 17'h0480a;
		 filter_in_data_log_force[ 763] <= 17'h180ab;
		 filter_in_data_log_force[ 764] <= 17'h05c45;
		 filter_in_data_log_force[ 765] <= 17'h007a8;
		 filter_in_data_log_force[ 766] <= 17'h19a08;
		 filter_in_data_log_force[ 767] <= 17'h07d32;
		 filter_in_data_log_force[ 768] <= 17'h1c20e;
		 filter_in_data_log_force[ 769] <= 17'h1d464;
		 filter_in_data_log_force[ 770] <= 17'h0772f;
		 filter_in_data_log_force[ 771] <= 17'h18e15;
		 filter_in_data_log_force[ 772] <= 17'h02019;
		 filter_in_data_log_force[ 773] <= 17'h046ee;
		 filter_in_data_log_force[ 774] <= 17'h1815b;
		 filter_in_data_log_force[ 775] <= 17'h062cb;
		 filter_in_data_log_force[ 776] <= 17'h1f99c;
		 filter_in_data_log_force[ 777] <= 17'h1a616;
		 filter_in_data_log_force[ 778] <= 17'h07fed;
		 filter_in_data_log_force[ 779] <= 17'h1ac27;
		 filter_in_data_log_force[ 780] <= 17'h1f287;
		 filter_in_data_log_force[ 781] <= 17'h06601;
		 filter_in_data_log_force[ 782] <= 17'h181be;
		 filter_in_data_log_force[ 783] <= 17'h047bf;
		 filter_in_data_log_force[ 784] <= 17'h01b05;
		 filter_in_data_log_force[ 785] <= 17'h1931b;
		 filter_in_data_log_force[ 786] <= 17'h07c13;
		 filter_in_data_log_force[ 787] <= 17'h1bff8;
		 filter_in_data_log_force[ 788] <= 17'h1dda4;
		 filter_in_data_log_force[ 789] <= 17'h06ff0;
		 filter_in_data_log_force[ 790] <= 17'h1851a;
		 filter_in_data_log_force[ 791] <= 17'h03d78;
		 filter_in_data_log_force[ 792] <= 17'h023b5;
		 filter_in_data_log_force[ 793] <= 17'h19022;
		 filter_in_data_log_force[ 794] <= 17'h07b5c;
		 filter_in_data_log_force[ 795] <= 17'h1bfb9;
		 filter_in_data_log_force[ 796] <= 17'h1e0e4;
		 filter_in_data_log_force[ 797] <= 17'h06cac;
		 filter_in_data_log_force[ 798] <= 17'h182c8;
		 filter_in_data_log_force[ 799] <= 17'h04837;
		 filter_in_data_log_force[ 800] <= 17'h01468;
		 filter_in_data_log_force[ 801] <= 17'h19a6c;
		 filter_in_data_log_force[ 802] <= 17'h07f5e;
		 filter_in_data_log_force[ 803] <= 17'h1ab83;
		 filter_in_data_log_force[ 804] <= 17'h1fc99;
		 filter_in_data_log_force[ 805] <= 17'h05935;
		 filter_in_data_log_force[ 806] <= 17'h18038;
		 filter_in_data_log_force[ 807] <= 17'h06382;
		 filter_in_data_log_force[ 808] <= 17'h1ec3b;
		 filter_in_data_log_force[ 809] <= 17'h1ba22;
		 filter_in_data_log_force[ 810] <= 17'h07b91;
		 filter_in_data_log_force[ 811] <= 17'h18d72;
		 filter_in_data_log_force[ 812] <= 17'h03010;
		 filter_in_data_log_force[ 813] <= 17'h02a25;
		 filter_in_data_log_force[ 814] <= 17'h190c9;
		 filter_in_data_log_force[ 815] <= 17'h07d89;
		 filter_in_data_log_force[ 816] <= 17'h1b13a;
		 filter_in_data_log_force[ 817] <= 17'h1fa2e;
		 filter_in_data_log_force[ 818] <= 17'h05754;
		 filter_in_data_log_force[ 819] <= 17'h180e2;
		 filter_in_data_log_force[ 820] <= 17'h06af2;
		 filter_in_data_log_force[ 821] <= 17'h1db11;
		 filter_in_data_log_force[ 822] <= 17'h1ce14;
		 filter_in_data_log_force[ 823] <= 17'h0718c;
		 filter_in_data_log_force[ 824] <= 17'h182bf;
		 filter_in_data_log_force[ 825] <= 17'h05063;
		 filter_in_data_log_force[ 826] <= 17'h0004a;
		 filter_in_data_log_force[ 827] <= 17'h1af76;
		 filter_in_data_log_force[ 828] <= 17'h07d0e;
		 filter_in_data_log_force[ 829] <= 17'h18d27;
		 filter_in_data_log_force[ 830] <= 17'h03703;
		 filter_in_data_log_force[ 831] <= 17'h01c2f;
		 filter_in_data_log_force[ 832] <= 17'h19ceb;
		 filter_in_data_log_force[ 833] <= 17'h07ff5;
		 filter_in_data_log_force[ 834] <= 17'h198b7;
		 filter_in_data_log_force[ 835] <= 17'h023f4;
		 filter_in_data_log_force[ 836] <= 17'h02dde;
		 filter_in_data_log_force[ 837] <= 17'h1934a;
		 filter_in_data_log_force[ 838] <= 17'h07f7e;
		 filter_in_data_log_force[ 839] <= 17'h1a0b9;
		 filter_in_data_log_force[ 840] <= 17'h0197b;
		 filter_in_data_log_force[ 841] <= 17'h03607;
		 filter_in_data_log_force[ 842] <= 17'h18fca;
		 filter_in_data_log_force[ 843] <= 17'h07ef3;
		 filter_in_data_log_force[ 844] <= 17'h1a2cf;
		 filter_in_data_log_force[ 845] <= 17'h01858;
		 filter_in_data_log_force[ 846] <= 17'h03555;
		 filter_in_data_log_force[ 847] <= 17'h1911c;
		 filter_in_data_log_force[ 848] <= 17'h07f75;
		 filter_in_data_log_force[ 849] <= 17'h19e73;
		 filter_in_data_log_force[ 850] <= 17'h0209a;
		 filter_in_data_log_force[ 851] <= 17'h02bb7;
		 filter_in_data_log_force[ 852] <= 17'h197c4;
		 filter_in_data_log_force[ 853] <= 17'h07ffa;
		 filter_in_data_log_force[ 854] <= 17'h194c8;
		 filter_in_data_log_force[ 855] <= 17'h031b9;
		 filter_in_data_log_force[ 856] <= 17'h0186f;
		 filter_in_data_log_force[ 857] <= 17'h1a5fa;
		 filter_in_data_log_force[ 858] <= 17'h07d4d;
		 filter_in_data_log_force[ 859] <= 17'h188f4;
		 filter_in_data_log_force[ 860] <= 17'h049ea;
		 filter_in_data_log_force[ 861] <= 17'h1faed;
		 filter_in_data_log_force[ 862] <= 17'h1beed;
		 filter_in_data_log_force[ 863] <= 17'h07243;
		 filter_in_data_log_force[ 864] <= 17'h180a2;
		 filter_in_data_log_force[ 865] <= 17'h064dc;
		 filter_in_data_log_force[ 866] <= 17'h1d485;
		 filter_in_data_log_force[ 867] <= 17'h1e527;
		 filter_in_data_log_force[ 868] <= 17'h058c2;
		 filter_in_data_log_force[ 869] <= 17'h18411;
		 filter_in_data_log_force[ 870] <= 17'h07a6d;
		 filter_in_data_log_force[ 871] <= 17'h1aac2;
		 filter_in_data_log_force[ 872] <= 17'h017a9;
		 filter_in_data_log_force[ 873] <= 17'h02c5d;
		 filter_in_data_log_force[ 874] <= 17'h19c79;
		 filter_in_data_log_force[ 875] <= 17'h07ea2;
		 filter_in_data_log_force[ 876] <= 17'h1895a;
		 filter_in_data_log_force[ 877] <= 17'h04e51;
		 filter_in_data_log_force[ 878] <= 17'h1eef4;
		 filter_in_data_log_force[ 879] <= 17'h1cf8d;
		 filter_in_data_log_force[ 880] <= 17'h064d2;
		 filter_in_data_log_force[ 881] <= 17'h18166;
		 filter_in_data_log_force[ 882] <= 17'h07795;
		 filter_in_data_log_force[ 883] <= 17'h1ade6;
		 filter_in_data_log_force[ 884] <= 17'h01820;
		 filter_in_data_log_force[ 885] <= 17'h0278d;
		 filter_in_data_log_force[ 886] <= 17'h1a2dd;
		 filter_in_data_log_force[ 887] <= 17'h07bc1;
		 filter_in_data_log_force[ 888] <= 17'h18390;
		 filter_in_data_log_force[ 889] <= 17'h05f8a;
		 filter_in_data_log_force[ 890] <= 17'h1d3a2;
		 filter_in_data_log_force[ 891] <= 17'h1ef30;
		 filter_in_data_log_force[ 892] <= 17'h049c9;
		 filter_in_data_log_force[ 893] <= 17'h18e46;
		 filter_in_data_log_force[ 894] <= 17'h08000;
		 filter_in_data_log_force[ 895] <= 17'h18e15;
		 filter_in_data_log_force[ 896] <= 17'h04b11;
		 filter_in_data_log_force[ 897] <= 17'h1ebba;
		 filter_in_data_log_force[ 898] <= 17'h1d97e;
		 filter_in_data_log_force[ 899] <= 17'h058d8;
		 filter_in_data_log_force[ 900] <= 17'h1878b;
		 filter_in_data_log_force[ 901] <= 17'h07f38;
		 filter_in_data_log_force[ 902] <= 17'h193c3;
		 filter_in_data_log_force[ 903] <= 17'h043ca;
		 filter_in_data_log_force[ 904] <= 17'h1f1bf;
		 filter_in_data_log_force[ 905] <= 17'h1d64a;
		 filter_in_data_log_force[ 906] <= 17'h05955;
		 filter_in_data_log_force[ 907] <= 17'h1883e;
		 filter_in_data_log_force[ 908] <= 17'h07fa7;
		 filter_in_data_log_force[ 909] <= 17'h18ffe;
		 filter_in_data_log_force[ 910] <= 17'h04c25;
		 filter_in_data_log_force[ 911] <= 17'h1e51d;
		 filter_in_data_log_force[ 912] <= 17'h1e536;
		 filter_in_data_log_force[ 913] <= 17'h04b71;
		 filter_in_data_log_force[ 914] <= 17'h1912d;
		 filter_in_data_log_force[ 915] <= 17'h07f38;
		 filter_in_data_log_force[ 916] <= 17'h185b6;
		 filter_in_data_log_force[ 917] <= 17'h0614c;
		 filter_in_data_log_force[ 918] <= 17'h1c747;
		 filter_in_data_log_force[ 919] <= 17'h00762;
		 filter_in_data_log_force[ 920] <= 17'h02ac5;
		 filter_in_data_log_force[ 921] <= 17'h1aa10;
		 filter_in_data_log_force[ 922] <= 17'h073ae;
		 filter_in_data_log_force[ 923] <= 17'h1802e;
		 filter_in_data_log_force[ 924] <= 17'h078f4;
		 filter_in_data_log_force[ 925] <= 17'h19f7e;
		 filter_in_data_log_force[ 926] <= 17'h03a65;
		 filter_in_data_log_force[ 927] <= 17'h1f3ae;
		 filter_in_data_log_force[ 928] <= 17'h1dce2;
		 filter_in_data_log_force[ 929] <= 17'h04d63;
		 filter_in_data_log_force[ 930] <= 17'h19319;
		 filter_in_data_log_force[ 931] <= 17'h07dbf;
		 filter_in_data_log_force[ 932] <= 17'h181f1;
		 filter_in_data_log_force[ 933] <= 17'h06e35;
		 filter_in_data_log_force[ 934] <= 17'h1af6b;
		 filter_in_data_log_force[ 935] <= 17'h02933;
		 filter_in_data_log_force[ 936] <= 17'h002e3;
		 filter_in_data_log_force[ 937] <= 17'h1d1bd;
		 filter_in_data_log_force[ 938] <= 17'h053d2;
		 filter_in_data_log_force[ 939] <= 17'h190a4;
		 filter_in_data_log_force[ 940] <= 17'h07dfe;
		 filter_in_data_log_force[ 941] <= 17'h18197;
		 filter_in_data_log_force[ 942] <= 17'h070f0;
		 filter_in_data_log_force[ 943] <= 17'h1a899;
		 filter_in_data_log_force[ 944] <= 17'h034d4;
		 filter_in_data_log_force[ 945] <= 17'h1f2ee;
		 filter_in_data_log_force[ 946] <= 17'h1e456;
		 filter_in_data_log_force[ 947] <= 17'h04142;
		 filter_in_data_log_force[ 948] <= 17'h19fe9;
		 filter_in_data_log_force[ 949] <= 17'h0755d;
		 filter_in_data_log_force[ 950] <= 17'h180ac;
		 filter_in_data_log_force[ 951] <= 17'h07d61;
		 filter_in_data_log_force[ 952] <= 17'h18ff6;
		 filter_in_data_log_force[ 953] <= 17'h058d4;
		 filter_in_data_log_force[ 954] <= 17'h1c5ee;
		 filter_in_data_log_force[ 955] <= 17'h016a5;
		 filter_in_data_log_force[ 956] <= 17'h00e55;
		 filter_in_data_log_force[ 957] <= 17'h1ce3e;
		 filter_in_data_log_force[ 958] <= 17'h050d0;
		 filter_in_data_log_force[ 959] <= 17'h196d4;
		 filter_in_data_log_force[ 960] <= 17'h07928;
		 filter_in_data_log_force[ 961] <= 17'h1802f;
		 filter_in_data_log_force[ 962] <= 17'h07cf5;
		 filter_in_data_log_force[ 963] <= 17'h18ee9;
		 filter_in_data_log_force[ 964] <= 17'h05d5a;
		 filter_in_data_log_force[ 965] <= 17'h1bca0;
		 filter_in_data_log_force[ 966] <= 17'h02524;
		 filter_in_data_log_force[ 967] <= 17'h1fb36;
		 filter_in_data_log_force[ 968] <= 17'h1e481;
		 filter_in_data_log_force[ 969] <= 17'h039ad;
		 filter_in_data_log_force[ 970] <= 17'h1ac0c;
		 filter_in_data_log_force[ 971] <= 17'h068e0;
		 filter_in_data_log_force[ 972] <= 17'h18899;
		 filter_in_data_log_force[ 973] <= 17'h07eed;
		 filter_in_data_log_force[ 974] <= 17'h180b8;
		 filter_in_data_log_force[ 975] <= 17'h078b7;
		 filter_in_data_log_force[ 976] <= 17'h19429;
		 filter_in_data_log_force[ 977] <= 17'h05992;
		 filter_in_data_log_force[ 978] <= 17'h1bcf6;
		 filter_in_data_log_force[ 979] <= 17'h02987;
		 filter_in_data_log_force[ 980] <= 17'h1f19f;
		 filter_in_data_log_force[ 981] <= 17'h1f2f0;
		 filter_in_data_log_force[ 982] <= 17'h0278a;
		 filter_in_data_log_force[ 983] <= 17'h1c016;
		 filter_in_data_log_force[ 984] <= 17'h0553a;
		 filter_in_data_log_force[ 985] <= 17'h19949;
		 filter_in_data_log_force[ 986] <= 17'h073d4;
		 filter_in_data_log_force[ 987] <= 17'h183c2;
		 filter_in_data_log_force[ 988] <= 17'h07fd8;
		 filter_in_data_log_force[ 989] <= 17'h18148;
		 filter_in_data_log_force[ 990] <= 17'h0791f;
		 filter_in_data_log_force[ 991] <= 17'h1908b;
		 filter_in_data_log_force[ 992] <= 17'h06240;
		 filter_in_data_log_force[ 993] <= 17'h1ade6;
		 filter_in_data_log_force[ 994] <= 17'h03fac;
		 filter_in_data_log_force[ 995] <= 17'h1d45a;
		 filter_in_data_log_force[ 996] <= 17'h016b4;
		 filter_in_data_log_force[ 997] <= 17'h1fe83;
		 filter_in_data_log_force[ 998] <= 17'h1ec9e;
		 filter_in_data_log_force[ 999] <= 17'h0275f;
		 filter_in_data_log_force[1000] <= 17'h1c5ff;
		 filter_in_data_log_force[1001] <= 17'h04ae2;
		 filter_in_data_log_force[1002] <= 17'h1a64c;
		 filter_in_data_log_force[1003] <= 17'h0663c;
		 filter_in_data_log_force[1004] <= 17'h18fad;
		 filter_in_data_log_force[1005] <= 17'h077e8;
		 filter_in_data_log_force[1006] <= 17'h18307;
		 filter_in_data_log_force[1007] <= 17'h07f94;
		 filter_in_data_log_force[1008] <= 17'h1802d;
		 filter_in_data_log_force[1009] <= 17'h07dde;
		 filter_in_data_log_force[1010] <= 17'h1861d;
		 filter_in_data_log_force[1011] <= 17'h07417;
		 filter_in_data_log_force[1012] <= 17'h1934e;
		 filter_in_data_log_force[1013] <= 17'h063f1;
		 filter_in_data_log_force[1014] <= 17'h1a5f0;
		 filter_in_data_log_force[1015] <= 17'h04f48;
		 filter_in_data_log_force[1016] <= 17'h1bc2c;
		 filter_in_data_log_force[1017] <= 17'h037e8;
		 filter_in_data_log_force[1018] <= 17'h1d448;
		 filter_in_data_log_force[1019] <= 17'h01f6f;
		 filter_in_data_log_force[1020] <= 17'h1ecca;
		 filter_in_data_log_force[1021] <= 17'h00732;
		 filter_in_data_log_force[1022] <= 17'h00481;
		 filter_in_data_log_force[1023] <= 17'h1f038;
		 filter_in_data_log_force[1024] <= 17'h01a8f;
		 filter_in_data_log_force[1025] <= 17'h1db3a;
		 filter_in_data_log_force[1026] <= 17'h02e61;
		 filter_in_data_log_force[1027] <= 17'h1c8a7;
		 filter_in_data_log_force[1028] <= 17'h03fa9;
		 filter_in_data_log_force[1029] <= 17'h1b8b1;
		 filter_in_data_log_force[1030] <= 17'h04e4d;
		 filter_in_data_log_force[1031] <= 17'h1ab5a;
		 filter_in_data_log_force[1032] <= 17'h00000;
		 filter_in_data_log_force[1033] <= 17'h00000;
		 filter_in_data_log_force[1034] <= 17'h00000;
		 filter_in_data_log_force[1035] <= 17'h00000;


        for (i = 0; i <= 1035; i = i + 1) begin
            input_data = filter_in_data_log_force[i][15:0];
            //#10;
				@(posedge clk);	
        end

        #100;
        $stop; 
    end

    // Monitor outputs
    initial begin
        $monitor("Time = %t, Input = %h, Output = %h, CE Out = %b",
                 $time, input_data, output_data, ce_out);
    end

endmodule
